`include "erasableMem.v"
`timescale 1 ns / 1 ps

module testmemReg ();
	reg clk;
	reg[2:0] bank;
	reg[9:0] memAddress;
	wire[16:0] dataOut;



endmodule // testmemReg