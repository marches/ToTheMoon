`timescale 1 ns / 1 ps

module memLogic (
	input[2:0] eBank,
	input[4:0] fBank,
	input superBank,
	input[11:0] memAddress,
	output[15:0] finalAddress	
);

endmodule