`timescale 1 ns / 1 ps

module erasableMem (
	input clk,    // Clock
	input[2:0] bank,
	input[9:0] memAddress,
	output[15:0] result	
);


endmodule